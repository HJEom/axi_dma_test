module sram #(parameter ADDR_WIDTH = 8, DATA_WIDTH = 8, DEPTH = 256) (
    input wire i_clk,
    input rstn,
    input ce,
    input wire [ADDR_WIDTH-1:0] i_addr, 
    input wire i_write,
    input wire [DATA_WIDTH-1:0] i_data,
    output reg [DATA_WIDTH-1:0] o_data 
    );

    (* ram_style = {"block"} *) reg [DATA_WIDTH-1:0] memory_array [0:DEPTH-1]; 

    always @ (posedge i_clk)
    begin
        if(ce) begin
        if(i_write) begin
            memory_array[i_addr] <= i_data;
            memory_array[i_addr+3] <= i_data;
        end
        else begin
            o_data <= memory_array[i_addr];
        end     
        end
    end
endmodule
